`ifdef DEFINES
`else
`define CLOCK_PERIOD 10  // DO NOT CHANGE
`define DEFINES 1
`define BITS 64
`define LOG_BITS 6
`endif
